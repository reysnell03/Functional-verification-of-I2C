class start_test extends test_base;

endclass
