package wb_pkg;
import ncsu_pkg::*;
`include"/mnt/ncsudrive/s/sreyya/745/project_2_provided_files/ece745_projects/proj_2/verification_ip/ncsu_pkg/ncsu_macros.svh"

`include "src/wb_configuration.svh"
`include "src/wb_transaction.svh"
`include "src/wb_driver.svh"
`include "src/wb_monitor.svh"
`include "src/wb_agent.svh"


endpackage
