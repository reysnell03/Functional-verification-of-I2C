class write_test extends test_base;

endclass
