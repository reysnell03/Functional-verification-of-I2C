class read_test extends test_base;

endclass
