class i2cmb_generator_test extends generator;
//`ncsu_register_object(i2cmb_generator_test)

endclass
